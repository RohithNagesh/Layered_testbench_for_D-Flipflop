interface intf(input bit clk);
  
  logic [2:0] D;
  logic reset;
  logic [2:0] Q;
  
endinterface